module CollisionDetection #(parameter N = 10)
			(reset, clk, pipe1_x, pipe1_y, pipe2_x, pipe2_y, pipe3_x, pipe3_y);
	input logic reset, clk;
	input logic [N-1 : 0] pipe1_x, pipe1_y0, pipe1_y1, 
								 pipe2_x, pipe2_y0, pipe2_y1,
								 pipe3_x, pipe3_y0, pipe3_y1;
	



endmodule
