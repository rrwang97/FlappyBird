module CollisionDetection();

endmodule 