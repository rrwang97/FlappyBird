module Randomizer();

endmodule 