module BirdDrawer();

endmodule 