module PipeDrawer();

endmodule 